
`include "rtl/design.sv"
`include "tb/top.sv"
